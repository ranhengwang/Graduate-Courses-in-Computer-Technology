`timescale 1ns/1ps

module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_size = 32;
reg [31:0] ROM_data[ROM_size-1:0];

always@(*)
	case(addr[8:2])	//Address Must Be Word Aligned.
		//LOOP3:
		//  addi $2, $0, 0x10
		0: data <= 32'b00100000000000100000000000010000;
		//  addi $3, $0, 0x0a
		1: data <= 32'b00100000000000110000000000001010;
		//  addi $7, $0, 0x0f
		2: data <= 32'b00100000000001110000000000001111;
		//  nop
		3: data <= 32'b00000000000000000000000000000000;
		//  nop
		4: data <= 32'b00000000000000000000000000000000;
		//  add $1, $2, $3
		5: data <= 32'b00000000010000110000100000100000;
		//  sub $4, $1, $3
		6: data <= 32'b00000000001000110010000000100010;
		//  and $6, $1, $7
		7: data <= 32'b00000000001001110011000000100100;
		//  addi $2, $0, 0x55
		8: data <= 32'b00100000000000100000000001010101;
		//  addi $3, $0, 0x10
		9: data <= 32'b00100000000000110000000000010000;
		//  addi $3, $0, 0x0a
		10: data <= 32'b00100000000000110000000000001010;
		//  addi $7, $0, 0x0f
		11: data <= 32'b00100000000001110000000000001111;
		//  addi $9, $0, 0x10
		12: data <= 32'b00100000000010010000000000010000;
		//  addi $11, $0, 0x11
		13: data <= 32'b00100000000010110000000000010001;
		//  nop
		14: data <= 32'b00000000000000000000000000000000;
		//  nop
		15: data <= 32'b00000000000000000000000000000000;
		//  add $1, $2, $3
		16: data <= 32'b00000000010000110000100000100000;
		//  sub $4, $1, $3
		17: data <= 32'b00000000001000110010000000100010;
		//  and $6, $1, $7
		18: data <= 32'b00000000001001110011000000100100;
		//  or $8, $1, $9
		19: data <= 32'b00000000001010010100000000100101;
		//  xor $10, $1, $11
		20: data <= 32'b00000000001010110101000000100110;
		//  addi $10, $0, 0x55AA
		21: data <= 32'b00100000000010100101010110101010;
		//  addi $2, $0, 0x20
		22: data <= 32'b00100000000000100000000000100000;
		//  addi $3, $0, 0x55
		23: data <= 32'b00100000000000110000000001010101;
		//  addi $9, $0, 0x00FF
		24: data <= 32'b00100000000010010000000011111111;
		//  sw $10, 0($2)
		25: data <= 32'b10101100010010100000000000000000;
		//  nop
		26: data <= 32'b00000000000000000000000000000000;
		//  nop
		27: data <= 32'b00000000000000000000000000000000;
		//  nop
		28: data <= 32'b00000000000000000000000000000000;
		//  lw $1, 0($2)
		29: data <= 32'b10001100010000010000000000000000;
		//  sub $7, $1, $3
		30: data <= 32'b00000000001000110011100000100010;
		//  and $6, $1, $7
		31: data <= 32'b00000000001001110011000000100100;
		//  or $8, $1, $9
		32: data <= 32'b00000000001010010100000000100101;
		//  addi $2, $0, 0x55
		33: data <= 32'b00100000000000100000000001010101;
		//  addi $4, $0, 0x0f
		34: data <= 32'b00100000000001000000000000001111;
		//  ori $3, $2, 0xaa
		35: data <= 32'b00110100010000110000000010101010;
		//  sub $5, $3, $4
		36: data <= 32'b00000000011001000010100000100010;
		//  nop
		37: data <= 32'b00000000000000000000000000000000;
		//  nop
		38: data <= 32'b00000000000000000000000000000000;
		//  addi $1, $0, 0xaa
		39: data <= 32'b00100000000000010000000010101010;
		//  addi $2, $0, 0x55
		40: data <= 32'b00100000000000100000000001010101;
		//  addi $4, $0, 0x0f
		41: data <= 32'b00100000000001000000000000001111;
		//  add $3, $2, $1
		42: data <= 32'b00000000010000010001100000100000;
		//  ori $6, $2, 1
		43: data <= 32'b00110100010001100000000000000001;
		//  sub $5, $3, $4
		44: data <= 32'b00000000011001000010100000100010;
		//  addi $1, $0, 0x55
		45: data <= 32'b00100000000000010000000001010101;
		//  addi $2, $0, 0xaa
		46: data <= 32'b00100000000000100000000010101010;
		//  addi $4, $0, 0x01
		47: data <= 32'b00100000000001000000000000000001;
		//  nop
		48: data <= 32'b00000000000000000000000000000000;
		//  sw $1, 0x08($0)
		49: data <= 32'b10101100000000010000000000001000;
		//  nop
		50: data <= 32'b00000000000000000000000000000000;
		//  nop
		51: data <= 32'b00000000000000000000000000000000;
		//  nop
		52: data <= 32'b00000000000000000000000000000000;
		//  lw $3, 0x08($0)
		53: data <= 32'b10001100000000110000000000001000;
		//  ori $6, $2, 0
		54: data <= 32'b00110100010001100000000000000000;
		//  sub $5, $3, $4
		55: data <= 32'b00000000011001000010100000100010;
		//  beq $3, $2, L1
		56: data <= 32'b00010000011000100000000000000000;
		//L1:
		//  add $4, $3, $2
		57: data <= 32'b00000000011000100010000000100000;
		//  sub $5, $3, $2
		58: data <= 32'b00000000011000100010100000100010;
		//  lw $1, 0($2)
		59: data <= 32'b10001100010000010000000000000000;
		//  sub $4, $1, $3
		60: data <= 32'b00000000001000110010000000100010;
		//  and $6, $1, $7
		61: data <= 32'b00000000001001110011000000100100;
		//  or $8, $1, $9
		62: data <= 32'b00000000001010010100000000100101;
		//  addi $1, $0, 0x89ABCDEF
		63: data <= 32'b001000000000000110001001101010111100110111101111;
		//  addi $2, $0, 0x12345678
		64: data <= 32'b001000000000001010010001101000101011001111000;
		//  sw $3, 8($0)
		65: data <= 32'b10101100000000110000000000001000;
		//  lw $4, 8($0)
		66: data <= 32'b10001100000001000000000000001000;
		//  nop
		67: data <= 32'b00000000000000000000000000000000;
		//  nop
		68: data <= 32'b00000000000000000000000000000000;
		//  nop
		69: data <= 32'b00000000000000000000000000000000;
		//  addi $7, $0, 0x20
		70: data <= 32'b00100000000001110000000000100000;
		//  addi $6, $0, 0x10
		71: data <= 32'b00100000000001100000000000010000;
		//  bne $6, $7, LOOP2
		72: data <= 32'b00010100110001110000000000000010;
		//  nop
		73: data <= 32'b00000000000000000000000000000000;
		//  nop
		74: data <= 32'b00000000000000000000000000000000;
		//LOOP2:
		//  beq $3, $4, LOOP3
		75: data <= 32'b00010000011001001111111110110100;
		//  nop
		76: data <= 32'b00000000000000000000000000000000;
		//  nop
		77: data <= 32'b00000000000000000000000000000000;
		//  nop
		78: data <= 32'b00000000000000000000000000000000;
		//LOOP1:
		//  j LOOP1
		79: data <= 32'b00001000000000000000000001001111;

	   default:	data <= 32'h8000_0000;
	endcase
endmodule
